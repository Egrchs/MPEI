// crc-16 x^16 + x^15 + x^2 + 1
module crc 
#(
    
) 
(
    input logic          CLK_I,
    input logic          RST_N_I,
    input logic [16 : 0] POLY_I
);
    
endmodule