`timescale 1ps/1ns

`define WAVES_FILE "dump/wave.vcd"

module tb();

endmodule