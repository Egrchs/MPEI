package fifo_sim_pkg;
    localparam real CLK_RD_PERIOD = 20;
    localparam real CLK_WR_PERIOD = 50;
endpackage