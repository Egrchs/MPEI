module dumpy(
    input  logic [7 : 0] data,
    output logic [7 : 0] data_o
);
    
endmodule