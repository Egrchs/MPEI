module qsubtract #(
                   parameter Q = 15,
                   parameter N = 32
                   )
  (
  input [N-1:0] a,
  input [N-1:0] b,
  output [N-1:0] c
  );

  reg [N-1:0] res;

  assign c = res;

  always @(a,b)
  begin
   // оба положительные или оба отрицательные
    if(a[N-1] == b[N-1])
    begin
      res[N-2:0] = a[N-2:0] - b[N-2:0];
      res[N-1] = a[N-1];
    end

   // один из операндов положительный
    else if(a[N-1] == 0 && b[N-1] == 1)
    begin
      if( a[N-2:0] > b[N-2:0] )
      begin
        res[N-2:0] = a[N-2:0] + b[N-2:0];
        res[N-1] = 1;
      end
      else
      begin
        res[N-2:0] = b[N-2:0] + a[N-2:0];
        if (res[N-2:0] == 0)
          res[N-1] = 0;
        else
          res[N-1] = 1;
        end
    end
    else
    begin
     if( a[N-2:0] > b[N-2:0] )
     begin
       res[N-2:0] = a[N-2:0] + b[N-2:0];
       if (res[N-2:0] == 0)
         res[N-1] = 0;
       else
         res[N-1] = 1;
       end
     else
     begin
       res[N-2:0] = b[N-2:0] + a[N-2:0];
       res[N-1] = 0;
     end
    end
  end
endmodule
