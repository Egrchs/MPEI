`include "cnt_FSM.v"

`timescale 1ns / 1ns

module tb_cnt_2_10_FSM();

reg iclk, irstn;
wire [7:0] oQ;

cnt_FSM DUT(.clk(iclk), .rst_n(irstn), .Q(oQ));

initial
begin
	iclk = 1'b0;
	irstn = 1'b1;
end

always #10 iclk = ~iclk;

initial
begin
	irstn = #20 ~irstn;
	irstn = #20 ~irstn;
end

initial
begin
	$dumpvars;
	#300 $finish;
end

endmodule
